
module procesamiento(







);



